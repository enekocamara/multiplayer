name=Multiplayer
port=12345
maxUsers=1000
queueSize=100
numOfRooms=3