name=Multiplayer
port=12346
maxUsers=1000
queueSize=100